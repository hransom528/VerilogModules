// XOR Gate

module xor(
	input x0, x1,
	output reg y);

	assign y = x0 ^ x1
endmodule